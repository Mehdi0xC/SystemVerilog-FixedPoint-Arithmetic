`ifndef _config_svh_
`define _config_svh_
`define F 17
`define N 32
`endif
