// Fixed-Point Testing Module for Multiplier with FixedPoint Size of N bits and Fraction Size of F bits
// Developed by Mehdi0xC, Winter 2018-2019
`include "config.svh"
module multiplier_test;
//##############################################################################################
//##############################################################################################
// PARAMETERs-----------------------------------------------------------------------------------
// INPUT AND OUTPUTS----------------------------------------------------------------------------
// VARIABLES -----------------------------------------------------------------------------------
	logic [31:0] a, b, c;
// MODULES INSTANTIATIONS-----------------------------------------------------------------------	
	multiplier  multiplier0 (
		.a(a), 
		.b(b), 
		.c(c)
	);
// INITIALIZATIONS------------------------------------------------------------------------------	
	initial
    begin								
		a[31:0] = 0;
        b[31:0] = 0;
        #100;
  	end
// MAIN-----------------------------------------------------------------------------------------
    always
    begin
        #100;
        a = 32'h0006487e;		
        b = 32'h00056fc2;
    end
//##############################################################################################
//##############################################################################################
endmodule
